* SPICE

V1 102 57 DC 10.0

R1 57 169 100
R2 170 102 100

.op
.tran 0 10ms 0ms 0.1ms
.end
