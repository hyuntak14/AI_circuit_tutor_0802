* SPICE

V1 168 115 DC 10.0

R1 115 111 100
R2 132 115 100
R3 121 118 100
V1 6 168 10.0

.op
.tran 0 10ms 0ms 0.1ms
.end
