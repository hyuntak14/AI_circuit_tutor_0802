* SPICE

V1 177 2 DC 10.0

R1 2 182 100
R2 182 115 100
R3 182 177 100
V1 2 177 10.0

.op
.tran 0 10ms 0ms 0.1ms
.end
