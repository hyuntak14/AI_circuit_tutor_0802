* SPICE

V1 4 4 DC 10.0

R1 4 4 100
R2 2 4 100

.op
.tran 0 10ms 0ms 0.1ms
.end
