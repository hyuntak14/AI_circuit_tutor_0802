* SPICE

V 0 0 DC 5


.op
.tran 0 10ms 0ms 0.1ms
.print 
.end
