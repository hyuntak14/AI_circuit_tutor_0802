* SPICE

V1 5 4 DC 10.0

R1 4 4 10
D2 4 2 Dmodel
R3 4 5 20

.op
.tran 0 10ms 0ms 0.1ms
.end
