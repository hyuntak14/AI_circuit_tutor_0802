* SPICE

V1 176 185 DC 5.0

R1 185 180 100
R2 180 176 100
R3 180 176 100
V1 184 176 5.0

.op
.tran 0 10ms 0ms 0.1ms
.end
