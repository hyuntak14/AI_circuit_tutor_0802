* SPICE

V1 176 443 DC 10.0

R1 443 180 100
R2 180 176 200
R3 180 176 300
V1 443 176 10.0

.op
.tran 0 10ms 0ms 0.1ms
.end
