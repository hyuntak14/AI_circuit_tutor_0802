* SPICE

V1 9 2 DC 10.0

R1 2 304 100
D2 304 9 Dmodel
D3 304 9 Dmodel
V1 2 9 10.0

.op
.tran 0 10ms 0ms 0.1ms
.end
