* SPICE

V1 175 443 DC 5.0

R1 443 180 100
R2 180 175 100
R3 180 175 100
V1 443 175 5.0

.op
.tran 0 10ms 0ms 0.1ms
.end
