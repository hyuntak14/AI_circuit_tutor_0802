* Multi-Power Circuit Netlist
* Generated with 1 power sources
* 
V1 185 9 5.0
R1 9 180 100.0
R2 180 185 100.0
R3 9 180 100.0
* 
.MODEL DMOD D
.MODEL LEDMOD D(IS=1E-12 N=2)
.END
