* Multi-Power Circuit Netlist
* Generated with 1 power sources
* Converted from: circuit5_superposition_a.graphml
* 
V1 1 2 15.0
R1 2 3 1000
R2 3 1 2000
R3 3 1 3000
* 
.MODEL DMOD D
.MODEL LEDMOD D(IS=1E-12 N=2)
.END