* Multi-Power Circuit Netlist
* Generated with 1 power sources
* 
V1 72 166 5.0
R1 72 166 100.0
R2 72 166 100.0
* 
.MODEL DMOD D
.MODEL LEDMOD D(IS=1E-12 N=2)
.END
