* SPICE

V1 102 177 DC 10.0

R1 177 171 100
R2 58 177 100
R3 171 102 100

.op
.tran 0 10ms 0ms 0.1ms
.end
