* SPICE

V1 102 177 DC 10.0

R1 177 170 1
D2 5 177 Dmodel
R3 163 102 2

.op
.tran 0 10ms 0ms 0.1ms
.end
