* SPICE

V1 177 187 DC 5.0

R1 187 182 100
R2 182 177 100
R3 178 182 100
V1 187 177 5.0

.op
.tran 0 10ms 0ms 0.1ms
.end
