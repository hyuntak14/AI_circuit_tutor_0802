* SPICE

V1 176 184 DC 5.0

L1 184 180 LEDmodel
C2 180 176 Cmodel
R3 180 176 100
V1 184 176 5.0

.op
.tran 0 10ms 0ms 0.1ms
.end
