* Multi-Power Circuit Netlist
* Generated with 3 power sources
* 
V1 2 4 0.2
V2 1 3 12.0
V3 2 6 12.0
R1 1 2 5100.0
R2 4 6 10000.0
X1 1 4 5 3 ua741
* 
.MODEL DMOD D
.MODEL LEDMOD D(IS=1E-12 N=2)
.END