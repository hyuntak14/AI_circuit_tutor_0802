* SPICE

V1 165 6 DC 5.6999999999999975

R1 6 114 100
R2 112 107 100
R3 112 107 100
V1 6 165 5.6999999999999975

.op
.tran 0 10ms 0ms 0.1ms
.end
