* Multi-Power Circuit Netlist
* Generated with 1 power sources
* Converted from: circuit3_Kirchhoff1.graphml
* 
V1 1 2 0.0
R1 2 3 1000
R2 3 1 2000
R3 3 1 3000
* 
.MODEL DMOD D
.MODEL LEDMOD D(IS=1E-12 N=2)
.END