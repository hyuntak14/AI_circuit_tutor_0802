* SPICE

V1 132 114 DC 10.0

R1 114 132 100
R2 113 132 20
R3 121 114 21
V1 122 132 10.0

.op
.tran 0 10ms 0ms 0.1ms
.end
