* Multi-Power Circuit Netlist
* Generated with 1 power sources
* Converted from: circuit6_oscilloscope.graphml
* 
V1 1 2 10.0
R1 2 1 3000
* 
.MODEL DMOD D
.MODEL LEDMOD D(IS=1E-12 N=2)
.END