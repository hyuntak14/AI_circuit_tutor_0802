* SPICE

V1 102 177 DC 10.0

R1 177 170 100
R2 5 177 100
R3 163 102 100

.op
.tran 0 10ms 0ms 0.1ms
.end
