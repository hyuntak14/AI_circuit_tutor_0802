* SPICE

V 4 2 DC 10.0

X2 5 2 10.0
X3 3 5 10.0
R4 4 3 100
R5 4 3 100

.op
.tran 0 10ms 0ms 0.1ms
.print v(1) v(2) v(3) 
.end
