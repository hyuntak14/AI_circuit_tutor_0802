* SPICE 

V 4 1 DC 10.0

L2 5 1 10
L3 3 5 10
R4 4 3 100
D5 3 4 10

.op
.tran 0 10ms 0ms 0.1ms
.print v(1) v(2) v(3) 
.end
