* SPICE

V1 156 6 DC 5.0

R1 6 114 50
R2 113 156 100
R3 113 156 200
V1 6 156 5.0

.op
.tran 0 10ms 0ms 0.1ms
.end
