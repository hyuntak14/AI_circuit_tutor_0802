* Multi-Power Circuit Netlist
* Generated with 1 power sources
* Converted from: circuit8_rectification.graphml
* 
V1 1 2 4.0
D1 2 3 DMOD
R1 3 1 2000
* 
.MODEL DMOD D
.MODEL LEDMOD D(IS=1E-12 N=2)
.END