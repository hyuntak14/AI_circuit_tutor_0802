* Multi-Power Circuit Netlist
* Generated with 1 power sources
* Converted from: circuit7_oscilloscope2.graphml
* 
V1 1 2 6.0
R1 2 3 1000
R2 3 1 2000
* 
.MODEL DMOD D
.MODEL LEDMOD D(IS=1E-12 N=2)
.END