* Multi-Power Circuit Netlist
* Generated with 1 power sources
* Converted from: circuit1_parellel_resistor.graphml
* 
V1 2 3 0.0
R1 3 2 2000
R2 3 2 3000
* 
.MODEL DMOD D
.MODEL LEDMOD D(IS=1E-12 N=2)
.END