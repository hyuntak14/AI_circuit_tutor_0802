* Multi-Power Circuit Netlist
* Generated with 1 power sources
* 
V1 6 167 5.0
R1 174 169 100.0
R2 6 174 100.0
R3 169 167 100.0
* 
.MODEL DMOD D
.MODEL LEDMOD D(IS=1E-12 N=2)
.END
