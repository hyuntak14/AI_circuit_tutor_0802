* Multi-Power Circuit Netlist
* Generated with 1 power sources
* Converted from: circuit2_series_resistor.graphml
* 
V1 2 3 0.0
R1 1 3 2.0
R2 1 2 2.0
* 
.MODEL DMOD D
.MODEL LEDMOD D(IS=1E-12 N=2)
.END