* SPICE

V1 162 196 DC 5.0

D1 196 162 Dmodel
R2 185 196 100
V1 185 162 5.0

.op
.tran 0 10ms 0ms 0.1ms
.end
