* SPICE 

V 4 5 DC 10.0


.op
.tran 0 10ms 0ms 0.1ms
.print 
.end
