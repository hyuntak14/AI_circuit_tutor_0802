* Multi-Power Circuit Netlist
* Generated with 1 power sources
* 
V1 2 3 6.0
R1 1 4 2000.0
R2 1 4 3000.0
* 
.MODEL DMOD D
.MODEL LEDMOD D(IS=1E-12 N=2)
.END